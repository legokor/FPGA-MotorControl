`timescale 1ns / 1ps

module test_pwm_generator();

// TODO

endmodule
